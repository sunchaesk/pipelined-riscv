
module pipeline_riscv_core (

                            );


endmodule
